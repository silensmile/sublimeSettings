always@(ways)
begin
	
end
function[:] name;
	
endfunction

if()
begin
	
end
else
begin
	
end
input[:] name;

output[:] name;

module name();
	
endmodule

reg[:] name;

